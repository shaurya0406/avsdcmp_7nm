** sch_path: /media/psf/avsdcmp_7nm/xschem/test/comparator_test.sch
**.subckt comparator_test
VDD VDD GND 0.7
VSS VSS GND 0
V1 Clk GND PULSE(0 0.7 10ps 5ps 5ps 240ps 500ps)
V2 Vin_p Vbias PULSE(-0.35 0.35 10ps 6000ps 10ps 10ps 6050ps)
V3 Vbias GND 0.35
V4 Vbias Vin_n PULSE(-0.35 0.35 10ps 6000ps 10ps 10ps 6050ps)
R1 Out_n VSS 10k m=1
R2 Out_p VSS 10k m=1
x1 VDD VSS Vin_p Out_n Vin_n Clk Out_p comparator
**** begin user architecture code


.control
run
TRAN 1p 6050p
plot Vin_p-Vin_n Out_p-Out_n Clk-4
plot Vin_p-Vin_n x1.pre_amp_p-x1.pre_amp_n Clk-4
.endc
.save all
.end


**** end user architecture code
**.ends

* expanding   symbol:  /media/psf/avsdcmp_7nm/xschem/src/comparator.sym # of pins=7
** sym_path: /media/psf/avsdcmp_7nm/xschem/src/comparator.sym
** sch_path: /media/psf/avsdcmp_7nm/xschem/src/comparator.sch
.subckt comparator VDD VSS Vin_p Out_n Vin_n Clk Out_p
*.iopin VDD
*.iopin VSS
*.ipin Vin_p
*.opin Out_n
*.ipin Vin_n
*.opin Out_p
*.ipin Clk
Xpfet1 Pre_Amp_n Clk_buf VDD VDD asap_7nm_pfet l=7e-009 nfin=7
Xpfet2 Pre_Amp_p Clk_buf VDD VDD asap_7nm_pfet l=7e-009 nfin=7
Xnfet1 Pre_Amp_n Vin_p net1 VSS asap_7nm_nfet l=7e-009 nfin=14
Xnfet2 Pre_Amp_p Vin_n net1 VSS asap_7nm_nfet l=7e-009 nfin=14
Xnfet3 net1 Clk_buf VSS VSS asap_7nm_nfet l=7e-009 nfin=14
Xpfet3 net2 net4 VDD VDD asap_7nm_pfet l=7e-009 nfin=2
Xpfet4 net3 net5 VDD VDD asap_7nm_pfet l=7e-009 nfin=2
Xpfet5 net5 Pre_Amp_n net2 VDD asap_7nm_pfet l=7e-009 nfin=4
Xpfet6 net4 Pre_Amp_p net3 VDD asap_7nm_pfet l=7e-009 nfin=4
Xnfet4 net5 Clk_n VSS VSS asap_7nm_nfet l=7e-009 nfin=10
Xnfet5 net5 net4 VSS VSS asap_7nm_nfet l=7e-009 nfin=10
Xnfet6 net4 net5 VSS VSS asap_7nm_nfet l=7e-009 nfin=10
Xnfet7 net4 Clk_n VSS VSS asap_7nm_nfet l=7e-009 nfin=10
Xpfet7 Clk_n Clk VDD VDD asap_7nm_pfet l=7e-009 nfin=14
Xnfet8 Clk_n Clk VSS VSS asap_7nm_nfet l=7e-009 nfin=14
x3 Out_p net6 VDD VSS buf8
x1 net6 net5 VDD VSS buf8
x2 Out_n net7 VDD VSS buf8
x10 net7 net4 VDD VSS buf8
x4 Clk_buf Clk VDD VSS buf8
.ends


* expanding   symbol:  buf8.sym # of pins=4
** sym_path: /media/psf/avsdcmp_7nm/xschem/lib/buf8.sym
** sch_path: /media/psf/avsdcmp_7nm/xschem/lib/buf8.sch
.subckt buf8 Out In VDD VSS
*.iopin VDD
*.iopin VSS
*.ipin In
*.opin Out
Xpfet1 net1 In VDD VDD asap_7nm_pfet l=7e-009 nfin=8
Xnfet1 net1 In VSS VSS asap_7nm_nfet l=7e-009 nfin=8
Xpfet2 Out net1 VDD VDD asap_7nm_pfet l=7e-009 nfin=8
Xnfet2 Out net1 VSS VSS asap_7nm_nfet l=7e-009 nfin=8
.ends

.GLOBAL GND
**** begin user architecture code

.subckt asap_7nm_pfet S G D B l=7e-009 nfin=8
	npmos_finfet S G D B BSIMCMG_osdi_P l=7e-009 nfin=8
.ends asap_7nm_pfet

.model BSIMCMG_osdi_P BSIMCMG_va (
+ TYPE = 0

************************************************************
*                         general                          *
************************************************************
+version = 107             bulkmod = 1               igcmod  = 1               igbmod  = 0
+gidlmod = 1               iimod   = 0               geomod  = 1               rdsmod  = 0
+rgatemod= 0               rgeomod = 0               shmod   = 0               nqsmod  = 0
+coremod = 0               cgeomod = 0               capmod  = 0               tnom    = 25
+eot     = 1e-009          eotbox  = 1.4e-007        eotacc  = 3e-010          tfin    = 6.5e-009
+toxp    = 2.1e-009        nbody   = 1e+022          phig    = 4.9278          epsrox  = 3.9
+epsrsub = 11.9            easub   = 4.05            ni0sub  = 1.1e+016        bg0sub  = 1.17
+nc0sub  = 2.86e+025       nsd     = 2e+026          ngate   = 0               nseg    = 5
+l       = 2.1e-008        xl      = 1e-009          lint    = -2.5e-009       dlc     = 0
+dlbin   = 0               hfin    = 3.2e-008        deltaw  = 0               deltawcv= 0
+sdterm  = 0               epsrsp  = 3.9             nfin    = 1
+toxg    = 1.8e-009
************************************************************
*                            dc                            *
************************************************************
+cit     = 0               cdsc    = 0.003469        cdscd   = 0.001486        dvt0    = 0.05
+dvt1    = 0.36            phin    = 0.05            eta0    = 0.094           dsub    = 0.24
+k1rsce  = 0               lpe0    = 0               dvtshift= 0               qmfactor= 0
+etaqm   = 0.54            qm0     = 2.183e-012      pqm     = 0.66            u0      = 0.0237
+etamob  = 4               up      = 0               ua      = 1.133           eu      = 0.05
+ud      = 0.0105          ucs     = 0.2672          rdswmin = 0               rdsw    = 200
+wr      = 1               rswmin  = 0               rdwmin  = 0               rshs    = 0
+rshd    = 0               vsat    = 60000           deltavsat= 0.17            ksativ  = 1.592
+mexp    = 2.491           ptwg    = 25              pclm    = 0.01            pclmg   = 1
+pdibl1  = 800             pdibl2  = 0.005704        drout   = 4.97            pvag    = 200
+fpitch  = 2.7e-008        rth0    = 0.15            cth0    = 1.243e-006      wth0    = 2.6e-007
+lcdscd  = 0               lcdscdr = 0               lrdsw   = 1.3             lvsat   = 1441
************************************************************
*                         leakage                          *
************************************************************
+aigc    = 0.007           bigc    = 0.0015          cigc    = 1               dlcigs  = 5e-009
+dlcigd  = 5e-009          aigs    = 0.006           aigd    = 0.006           bigs    = 0.001944
+bigd    = 0.001944        cigs    = 1               cigd    = 1               poxedge = 1.152
+agidl   = 2e-012          agisl   = 2e-012          bgidl   = 1.5e+008        bgisl   = 1.5e+008
+egidl   = 1.142           egisl   = 1.142
************************************************************
*                            rf                            *
************************************************************
************************************************************
*                         junction                         *
************************************************************
************************************************************
*                       capacitance                        *
************************************************************
+cfs     = 0               cfd     = 0               cgso    = 1.6e-010        cgdo    = 1.6e-010
+cgsl    = 0               cgdl    = 0               ckappas = 0.6             ckappad = 0.6
+cgbo    = 0               cgbl    = 0
************************************************************
*                       temperature                        *
************************************************************
+tbgasub = 0.000473        tbgbsub = 636             kt1     = 0               kt1l    = 0
+ute     = -1.2            utl     = 0               ua1     = 0.001032        ud1     = 0
+ucste   = -0.004775       at      = 0.001           ptwgt   = 0.004           tmexp   = 0
+prt     = 0               tgidl   = -0.007          igt     = 2.5
************************************************************
*                          noise                           *
************************************************************
**)
.control
pre_osdi ~/ASAP7_FinFET_Inverter_Characterization/Xschem_ASAP7/bsimcmg_arch64.osdi
.endc



.subckt asap_7nm_nfet S G D B l=7e-009 nfin=8
	nnmos_finfet S G D B BSIMCMG_osdi_N l=7e-009 nfin=8
.ends asap_7nm_nfet

.model BSIMCMG_osdi_N BSIMCMG_va (
+ TYPE = 1
************************************************************
*                         general                          *
************************************************************
+version = 107             bulkmod = 1               igcmod  = 1               igbmod  = 0
+gidlmod = 1               iimod   = 0               geomod  = 1               rdsmod  = 0
+rgatemod= 0               rgeomod = 0               shmod   = 0               nqsmod  = 0
+coremod = 0               cgeomod = 0               capmod  = 0               tnom    = 25
+eot     = 1e-009          eotbox  = 1.4e-007        eotacc  = 1e-010          tfin    = 6.5e-009
+toxp    = 2.1e-009        nbody   = 1e+022          phig    = 4.2466          epsrox  = 3.9
+epsrsub = 11.9            easub   = 4.05            ni0sub  = 1.1e+016        bg0sub  = 1.17
+nc0sub  = 2.86e+025       nsd     = 2e+026          ngate   = 0               nseg    = 5
+l       = 2.1e-008        xl      = 1e-009          lint    = -2e-009         dlc     = 0
+dlbin   = 0               hfin    = 3.2e-008        deltaw  = 0               deltawcv= 0
+sdterm  = 0               epsrsp  = 3.9             nfin    = 1
+toxg    = 1.80e-009
************************************************************
*                            dc                            *
************************************************************
+cit     = 0               cdsc    = 0.01            cdscd   = 0.01            dvt0    = 0.05
+dvt1    = 0.47            phin    = 0.05            eta0    = 0.07            dsub    = 0.35
+k1rsce  = 0               lpe0    = 0               dvtshift= 0               qmfactor= 2.5
+etaqm   = 0.54            qm0     = 0.001           pqm     = 0.66            u0      = 0.0303
+etamob  = 2               up      = 0               ua      = 0.55            eu      = 1.2
+ud      = 0               ucs     = 1               rdswmin = 0               rdsw    = 200
+wr      = 1               rswmin  = 0               rdwmin  = 0               rshs    = 0
+rshd    = 0               vsat    = 70000           deltavsat= 0.2             ksativ  = 2
+mexp    = 4               ptwg    = 30              pclm    = 0.05            pclmg   = 0
+pdibl1  = 0               pdibl2  = 0.002           drout   = 1               pvag    = 0
+fpitch  = 2.7e-008        rth0    = 0.225           cth0    = 1.243e-006      wth0    = 2.6e-007
+lcdscd  = 5e-005          lcdscdr = 5e-005          lrdsw   = 0.2             lvsat   = 0
************************************************************
*                         leakage                          *
************************************************************
+aigc    = 0.014           bigc    = 0.005           cigc    = 0.25            dlcigs  = 1e-009
+dlcigd  = 1e-009          aigs    = 0.0115          aigd    = 0.0115          bigs    = 0.00332
+bigd    = 0.00332         cigs    = 0.35            cigd    = 0.35            poxedge = 1.1
+agidl   = 1e-012          agisl   = 1e-012          bgidl   = 10000000        bgisl   = 10000000
+egidl   = 0.35            egisl   = 0.35
************************************************************
*                            rf                            *
************************************************************
************************************************************
*                         junction                         *
************************************************************
************************************************************
*                       capacitance                        *
************************************************************
+cfs     = 0               cfd     = 0               cgso    = 1.6e-010        cgdo    = 1.6e-010
+cgsl    = 0               cgdl    = 0               ckappas = 0.6             ckappad = 0.6
+cgbo    = 0               cgbl    = 0
************************************************************
*                       temperature                        *
************************************************************
+tbgasub = 0.000473        tbgbsub = 636             kt1     = 0               kt1l    = 0
+ute     = -0.7            utl     = 0               ua1     = 0.001032        ud1     = 0
+ucste   = -0.004775       at      = 0.001           ptwgt   = 0.004           tmexp   = 0
+prt     = 0               tgidl   = -0.007          igt     = 2.5
************************************************************
*                          noise                           *
************************************************************
**)
.control
pre_osdi ~/ASAP7_FinFET_Inverter_Characterization/Xschem_ASAP7/bsimcmg_arch64.osdi
.endc


**** end user architecture code
.end
